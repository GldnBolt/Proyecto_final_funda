module top(
    input  logic        clk,
    input  logic        reset,
    output logic [31:0] WriteData,
    output logic [31:0] DataAdr,
    output logic        MemWrite,
	 
	     // --- Salidas VGA ---
    output vgaclk,
    output hsync,
    output vsync,
    output sync_b,
    output blank_b,
    output [7:0] r, // << Salidas finales multiplexadas
    output [7:0] g,
    output [7:0] b
	 
);


    // Señales internas
    logic [31:0] PC, Instr, ReadData;

    // Señal interna para el contador de ciclos
    logic [7:0] cycle_counter;  // Instancia de un contador de 8 bits (puedes ajustarlo a más bits si necesitas más capacidad)
	 
	 // --- Señales Internas ---
    wire [9:0] x, y; // Coordenadas desde vgaController



    // --- Señales RGB intermedias para los dos generadores de video ---
	 wire [7:0] start_r, start_g, start_b; // RGB desde startScreen


    // --- Instancia PLL (Sin cambios) ---
    pll vgapll(.inclk0(clk), .c0(vgaclk));

    // --- Instancia Controlador VGA (Sin cambios) ---
    // Genera vgaclk, hsync, vsync, sync_b, blank_b, x, y
    vgaController vgaCont(
        .vgaclk(vgaclk), .hsync(hsync), .vsync(vsync), .sync_b(sync_b),
        .blank_b(blank_b), .x(x), .y(y)
    );
	 
	 startScreen initialScreenDrawer (
        .x(x),                         // Coordenada X desde vgaController
        .y(y),                         // Coordenada Y desde vgaController
        .visible(1), // Se muestra solo si la FSM está en P_INICIO
        .r(start_r),                   // Salida R de la pantalla de inicio
        .g(start_g),                   // Salida G de la pantalla de inicio
        .b(start_b)                    // Salida B de la pantalla de inicio
    );

    // --- Multiplexor de Salida RGB Final ---
    // Si es el estado inicial, usa los colores de startScreen, si no, los de videoGen (juego)
    assign r = start_r ;
    assign g = start_g ;
    assign b = start_b ;


    // Instancia del procesador
    arm arm0 (
        .clk       (clk),
        .reset     (reset),
        .PC        (PC),
        .Instr     (Instr),
        .MemWrite  (MemWrite),
        .ALUResult (DataAdr),
        .WriteData (WriteData),
        .ReadData  (ReadData)
    );

    // Memoria de instrucciones (imem.sv)
    // Asegúrate de que en imem.sv tengas:
    //   initial $readmemh("ROM.dat", RAM);
	     imem imem0 (
        .a  (PC),    // byte-address de instrucción
        .rd (Instr)  // instrucción de 32 bits
    );

    // Memoria de datos (dmem.sv)
    // Memoria de datos de dos puertos (dmem.sv)
    dmem dmem0 (
        .clk    (clk),        // reloj
        .we     (MemWrite),   // habilita escritura en puerto 0
        .addr0  (DataAdr),    // dirección byte-address puerto 0
        .wd0    (WriteData),  // dato a escribir            puerto 0
        .rd0    (ReadData),   // dato leído                 puerto 0

        .addr1  (32'b0),      // puerto 1 sólo lectura: dirección fija a 0
        .rd1    ()            // puerto 1 sólo lectura: salida no conectada
    );


endmodule
